module mux4in (x, sel, y);
    input [3:0] x;                      // sel selects the exit (x[3], x[2], x[1], x[0]).
    input [1:0] sel;
    output reg y;

    reg curr;                           // Curr is the register the mux is copying currently.

    always @(sel or x) begin
        if (sel == 0)
            assign y = x[0];
        else if (sel == 1)
            assign y = x[1];
        else if (sel == 2)
            assign y = x[2];
        else if (sel == 3)
            assign y = x[3];

    end

endmodule