module decoder4out(x1, x2, y1, y2, y3, y4);
    input x1, x2;
    output y1, y2, y3, y4;

endmodule